module hello;
    initial begin
        $display("hello world");
        $finish;
    end
endmodule  
