module test (a,b,c,d,e);  
input[3:0]a,b,c;
output[3:0]d,e;
wire[3:0]a,b,c,d,e;
endmodule
